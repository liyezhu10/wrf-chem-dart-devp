netcdf simple{

dimensions:
lat   = 4;
lon   = 2;
time = UNLIMITED ; //(1 currently)
variables:

double temp(time,lon,lat);
temp:units = "palm trees" ;
temp:long_name = "ambient spectacular temperature from some really great planet and season" ;
temp:short_name = "temperature" ;

float time(time);
time:units = "hours" ;

//global attributes:

:title = "simple_file" ;

data:
time = 1 ;

temp = 
   1.0, 2.0, 3.0,  4.0,  
   5.0, 6.0, 7.0,  8.0;

}
